----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 29.04.2017 18:34:01
-- Design Name: 
-- Module Name: player1_rom - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SilverSurfer_fire_rom is
    Port ( address : in STD_LOGIC_VECTOR (9 downto 0);
           pixel_out : out STD_LOGIC_VECTOR (11 downto 0));
end SilverSurfer_fire_rom;

architecture Behavioral of SilverSurfer_fire_rom is

type row_type is array(0 to 19) of std_logic_vector(11 downto 0);
type SilverSurfer_fire_rom_type is array(0 to 19) of row_type;
signal row : row_type;

constant SilverSurfer_fire_ROM : SilverSurfer_fire_rom_type := 
(
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "110011011110", "101111101111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011010111101", "001110111101", "001011011111", "101111101111", "110011011110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "001111001110", "001111011111", "001111101111", "001111111111", "001011011111", "001110111101", "011110111101", "110111011101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111011111110", "001111001110", "001111111111", "011111111111", "011111111111", "010011111111", "001111111111", "001111101111", "001111101111", "010011011110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "011010111110", "001111101111", "011011111111", "010011111111", "011111111111", "111011111111", "010011111111", "011111111111", "011111111111", "001111111111", "001111001110", "111011101110", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111011111111", "011011011110", "001111101111", "100011111111", "011111111111", "111111111111", "111111111111", "111011111111", "011111111111", "010011111111", "011011111111", "001111101111", "010110101101", "111111111110", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "101111101111", "010011101111", "001111111111", "010011111111", "111011111111", "111111111111", "111111111111", "111111111111", "111111111111", "100011111111", "100011111111", "001111101111", "010011001110", "110011011110", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "101011101111", "001011011111", "001111111111", "010011111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011111111", "010011111111", "001111111111", "001011011111", "100111011110", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "101111011110", "001110111110", "001111101111", "011011111111", "011111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010111111111", "001111111111", "001011101111", "101011101111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111011011110", "010110011100", "001111101111", "100011111111", "010111111111", "100011111111", "111011111111", "111111111111", "111111111111", "100011111111", "011011111111", "001111101111", "001111001110", "101111011110", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "110011011101", "001111001110", "001111111111", "011111111111", "011111111111", "010111111111", "111011111111", "100011111111", "010111111111", "100011111111", "001111101111", "011010111110", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "010111011111", "001111101111", "001111101111", "001111111111", "010111111111", "011111111111", "011111111111", "001111111111", "010011011110", "110111011101", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011111111", "011010111110", "001111001110", "001011101111", "001111111111", "001111101111", "001111101111", "001011001110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "101011001110", "100111101111", "001011101111", "001111001110", "010110111110", "110111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100111101111", "101111011110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111")

);

begin

row <= SilverSurfer_fire_ROM(conv_integer(address(9 downto 5)));
pixel_out <= row(conv_integer(address(4 downto 0)));

end Behavioral;