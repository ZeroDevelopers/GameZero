----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 29.04.2017 18:34:01
-- Design Name: 
-- Module Name: player1_rom - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity GreenGoblin_rom is
    Port ( address : in STD_LOGIC_VECTOR (11 downto 0);
           pixel_out : out STD_LOGIC_VECTOR (11 downto 0));
end GreenGoblin_rom;

architecture Behavioral of GreenGoblin_rom is

type row_type is array(0 to 63) of std_logic_vector(11 downto 0);
type GreenGoblin_rom_type is array(0 to 63) of row_type;
signal row : row_type;

constant GREENGOBLIN_ROM : GreenGoblin_rom_type := 
(
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "111111111111", "011101110111", "010101010101", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "011000011001", "010001000100", "011000011001", "100000111100", "001000100010", "001111001010", "001000100010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "001100000111", "010100001001", "100000111100", "100000111100", "010100001001", "001000100010", "001111001010", "001000100010", "100000111100", "011000011001", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "010100001001", "000110010101", "010100001001", "010100001001", "001000100010", "000110010101", "001111001010", "001000100010", "100000111100", "010100001001", "011000011001", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011000011001", "000110010101", "001111001010", "001000000110", "001000000110", "001000100010", "001111001010", "001111001010", "001000100010", "010100001001", "100000111100", "100000111100", "010100001001", "001100000111", "010001000100", "111111111111", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "010100001001", "111011101110", "000110010101", "000001100011", "001000000110", "000001100011", "001111001010", "001111001010", "001000100010", "001000100010", "001000100010", "100000111100", "100000111100", "010100001001", "001000000110", "001000000011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "001000100010", "001000100010", "000110010101", "000001000010", "111011101110", "001000000110", "000110010101", "001111001010", "000110010101", "001000100010", "010100001001", "001000000110", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000000110", "010100001001", "100000111100", "100101001101", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "000110010110", "001000100010", "111011101110", "001111001010", "111011101110", "111011101110", "010100001001", "001111001010", "001111001010", "000001100011", "001000100010", "100000111100", "010100001001", "001000000110", "001000100010", "000001100011", "000001100011", "000001000010", "001000100010", "001000100010", "001000000110", "100000111100", "100000111100", "011000011001", "011001100110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110011011011", "010001000100", "001111001010", "001000100010", "000110010101", "001111001010", "000110010101", "000001100011", "001111001010", "000110010101", "001111001010", "000001000010", "001000100010", "100000111100", "100000111100", "010100001001", "001000100010", "001111001010", "001111001010", "000110010101", "000001000010", "000001000010", "001000100010", "010001000100", "010001000100", "100101001101", "011000101010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "010001000100", "001000100010", "001111001010", "000001100011", "001000100010", "000001100011", "000110010101", "000001100011", "000110010101", "001000100010", "000110010101", "001000100010", "010100001001", "010100001001", "010100001001", "001000100010", "000110010101", "001111001010", "001111001010", "000110010101", "000001100011", "000001000010", "001100110011", "101111001001", "101111001001", "010101010101", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "000110010110", "001111001010", "001000100010", "000110010101", "000001100011", "001000100010", "001111001010", "000001100011", "000001000010", "000110010101", "000001000010", "001000100010", "001000000110", "010100001001", "001000000110", "000100000011", "001000100010", "000001100011", "000110010101", "000110010101", "000001100011", "000001100011", "001000100010", "000101000010", "001101100100", "010101010101", "101111001001", "111011101100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "000101000010", "000001100011", "000110010101", "001000100010", "000001000010", "000001100011", "001000100010", "000110010101", "001000100010", "001000100010", "000001000010", "000001000010", "001000100010", "001000000110", "001000000110", "010100001001", "001000000110", "001000100010", "000001000010", "000001100011", "000001100011", "000001100011", "001000100010", "000001000010", "000001100011", "001111001010", "000101100011", "001101100100", "100010001000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "001111011011", "000001100011", "001111001010", "001111001010", "000110010101", "001000100010", "000001000010", "001000100010", "001000100010", "000001001001", "001000100010", "001000100010", "001000000110", "010100001001", "100000111100", "100000111100", "100000111100", "001000000110", "001000100010", "000001000010", "001000100010", "001000100010", "001000100010", "000001000010", "000001000010", "000001000010", "000001100011", "000110010101", "000001000010", "000101000010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "000110010101", "000001100011", "001111001010", "000110010101", "000001100011", "000101000010", "001100110011", "001000100010", "001000000110", "001000100010", "000001001001", "001000100010", "001000100010", "001000000110", "010100001001", "100000111100", "100000111100", "001000000110", "000100000011", "001000100010", "000001000010", "000001000010", "000110010101", "000110010101", "000110010101", "000001100011", "000001000010", "000001100011", "000001000010", "000001100011", "000001100011", "001111011011", "111111111111", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "000101100011", "000110010101", "000001000010", "000001100011", "000001100011", "000101000010", "011001100110", "110011011010", "011001100110", "001100000111", "100000111100", "001000100010", "000001001001", "000001001001", "001000100010", "001000100010", "010100001001", "010100001001", "010100001001", "000100000011", "000100000011", "001000100010", "001000100010", "000001100011", "001111001010", "001111001010", "000110010101", "000001100011", "001000100010", "000001100011", "000001000010", "000110010101", "000001100011", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "000001000010", "000110010101", "001111001010", "000110010101", "001000100010", "011001100110", "110111101100", "111111111110", "110111101100", "011001100110", "001100000111", "100000111100", "001000100010", "001000100010", "000001001001", "000001001001", "001000100010", "001000100010", "001000000110", "001000000110", "000100000011", "000100000011", "000100000011", "001000100010", "000001000010", "001111001010", "001111001010", "000001100011", "001000100010", "000001000010", "000110010101", "001111001010", "000110010101", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "001000100010", "000001100011", "001111001010", "000101100011", "011001100110", "110111101100", "111111111111", "111111111111", "111111111111", "110111101100", "011101110111", "010100001001", "010100001001", "000100000011", "001000100010", "001000100010", "000001001001", "000001001001", "001000100010", "001000100010", "001000100010", "001000000110", "001000000110", "000100000011", "001000100010", "000001000010", "000001000010", "000001000010", "001000100010", "000110010101", "001111001010", "001111001010", "000110010101", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "100101001101", "100000111100", "001000100010", "000110010110", "011001100110", "110111101100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010000110101", "001100000111", "001000000110", "000100000011", "000100000011", "001000100010", "001000100010", "000001001001", "000001001001", "000001001001", "001000100010", "001000100010", "000100000011", "100010100100", "001000100010", "001000100010", "001000100010", "001000100010", "000110010101", "001000100010", "001000100010", "001000100010", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "010100001001", "000100000011", "100000111100", "010001000100", "110111101011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "001000000011", "010100001001", "010100001001", "100000111100", "010100001001", "001000100010", "001000100010", "001000100010", "000001001001", "000001001001", "001000100010", "001000100010", "100010100100", "100010100100", "100010100100", "001000100010", "001000100010", "100000111100", "010100001001", "001000000110", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "001000000110", "010100001001", "000100000011", "010101010101", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101100", "010001000100", "001000100010", "001000100010", "001000100010", "001000100010", "000100000011", "000001001001", "000010001110", "001000100010", "001000100010", "000001001001", "000001001001", "001000100010", "001000100010", "001000100010", "100000111100", "100000111100", "001000000110", "000100000011", "001000000011", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "001000100010", "100000111100", "001000000110", "010001000100", "110111101011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "000001001001", "000010001110", "000010001110", "000010001110", "000010001110", "000010001110", "000001001001", "000100000011", "001000100010", "001000100010", "001000100010", "000001001001", "000001001001", "001000100010", "001000000110", "100000111100", "010100001001", "001000000110", "001100110011", "110011011001", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "100000111100", "100000111100", "100000111100", "100101001101", "011001100110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "001000100010", "000001001001", "000010001110", "000010001110", "000001001001", "001000100010", "001000100010", "001000100010", "010100001001", "001000100010", "100010100100", "001000100010", "001000100010", "001000100010", "001000100010", "100000111100", "100000111100", "000100000011", "001000100010", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "100000111100", "001000000110", "001000000110", "001000000110", "100101001101", "100010001000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "111111111111", "110111101100", "010001000100", "010100001001", "001000100010", "001000100010", "001000100010", "001000100010", "010100001001", "100000111100", "100000111100", "010100001001", "001000100010", "100010100100", "100010100100", "001000100010", "001000000110", "010100001001", "100000111100", "001000000110", "000100000011", "001000100010", "001000100010", "001000100010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "100101001101", "001000000110", "001100000111", "010001000100", "010101010101", "011101110111", "110111101011", "111111111111", "111111111111", "100110011001", "011001100110", "010101010101", "010101010101", "111111111111", "011001100110", "100101001101", "010100001001", "100000111100", "100000111100", "100000111100", "100000111100", "010100001001", "010100001001", "001000100010", "001000100010", "000001100011", "001000100010", "001000100010", "100000111100", "100000111100", "100000111100", "100000111100", "010100001001", "001000100010", "001000100010", "000001001001", "001000100010", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "100000111100", "001000000110", "010001000100", "110011011011", "110111101100", "110111011011", "110011011011", "011101110111", "010001000100", "000101100011", "000110010101", "001111001010", "001111001010", "010001000100", "001000100010", "001000100010", "100000111100", "001000000110", "000100000011", "000100000011", "001000000110", "100000111100", "001000100010", "000110010101", "001111001010", "001111001010", "001000100010", "100000111100", "001000100010", "010100001001", "100000111100", "100000111100", "010100001001", "001000100010", "001000100010", "000001001001", "001000100010", "001000100010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "100101001101", "001000000110", "010001000100", "110011011011", "110111101011", "011101110111", "010001000100", "000101100011", "000110010101", "001111001010", "001111001010", "001111001010", "000110010101", "001111001010", "000110010101", "000001000010", "001000100010", "010100001001", "001000000110", "001000000110", "100000111100", "001000100010", "000001100011", "000001100011", "001111001010", "000110010101", "000001100011", "001000100010", "001000100010", "100000111100", "100000111100", "010100001001", "010100001001", "001000100010", "001000100010", "000001001001", "000001001001", "001000100010", "111111111111", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "100101001101", "001000100010", "010001000100", "001101100100", "000101100011", "000001000010", "000001000010", "000001100011", "000001100011", "000001100011", "000001000010", "000001000010", "000001100011", "000001000010", "000001100011", "001000100010", "001000000110", "010100001001", "010100001001", "001000100010", "000001100011", "000110010101", "000001000010", "000001000010", "000001100011", "000001100011", "001000100010", "100000111100", "001000100010", "100000111100", "001000100010", "010100001001", "001000100010", "000001001001", "001000100010", "000001001001", "001100110011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "001000100010", "001111001010", "001111001010", "000110010101", "000001100011", "000001100011", "000001000010", "000001000010", "000001000010", "000001100011", "000110010101", "000001000010", "000001100011", "000110010101", "000001100011", "001000100010", "001000000110", "001000000110", "001000100010", "000110010101", "001111001010", "000110010101", "000001000010", "000001000010", "000001100011", "001111001010", "001000100010", "100000111100", "001000100010", "010100001001", "001000100010", "000001001001", "000001001001", "001000100010", "000001001001", "000001001010", "111111111111", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "001111001010", "000110010101", "000001100011", "000001100011", "000110010101", "000110010101", "001111001010", "001111001010", "001111001010", "001111001010", "000001100011", "000110010101", "001111001010", "000001000010", "001000100010", "001000000110", "001000000110", "001000100010", "000001100011", "001111001010", "000001100011", "001111001010", "001111001010", "000001000010", "000110010101", "000001100011", "001000100010", "001000100010", "001000100010", "000001001001", "000001001001", "000001001001", "000001001001", "001000100010", "000001001001", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "000110010101", "000001100011", "000001000010", "000001000010", "000001100011", "000001100011", "000110010101", "001111001010", "001111001010", "000110010101", "000110010101", "000001100011", "000001000010", "000001000010", "001000100010", "001000000110", "001000000110", "001000100010", "000001000010", "000001100011", "000001100011", "001111001010", "000110010101", "000001000010", "000001100011", "000001000010", "000001000010", "001000100010", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "001000100010", "000001001001", "000001001010", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000101000010", "000001000010", "000001000010", "001000100010", "000001000010", "000001000010", "000001000010", "000001100011", "000001100011", "000001100011", "000001100011", "000001100011", "000001000010", "000001100011", "001000100010", "000100000011", "000100000011", "001000100010", "000001000010", "000001000010", "000001000010", "000110010101", "000110010101", "000001000010", "000001000010", "000001000010", "001000100010", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "001000100010", "000001001010", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "001000100010", "000001000010", "000001000010", "001000100010", "001000100010", "001000100010", "000001000010", "000001000010", "000001000010", "000001100011", "000001000010", "000001100011", "001000100010", "010000110101", "010101010101", "010101010101", "010000110101", "001000100010", "000001000010", "000110010101", "001000100010", "001000100010", "000001000010", "000001000010", "001000100010", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "000001001010", "010001000100", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "000101000010", "000001100011", "000001000010", "000001100011", "000001000010", "001000100010", "001000100010", "010001000100", "010101010101", "000101000010", "010001000100", "010101010101", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "001000100010", "000001100011", "000001000010", "001000100010", "000001000010", "000001000010", "001000100010", "000001001001", "000001001001", "000001001001", "000001001001", "000001001001", "000001001010", "010001000100", "011101110111", "110111101011", "111011111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "000001100011", "000001000010", "000110010101", "001111001010", "000001000010", "010001000100", "110011011011", "111111111111", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001100110", "000101000010", "000001000010", "000001000010", "000001000010", "000110010101", "000001100011", "001000100010", "000001001001", "000001001001", "000001001010", "010001000100", "011101110111", "110111101011", "111011111101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000101000010", "000001100011", "000110010101", "001111001010", "001111001010", "010001000100", "110111101100", "111111111111", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101100", "010001000100", "000001000010", "000001100011", "000001000010", "001111001010", "000110010101", "000001000010", "001000100010", "010001000100", "011101110111", "110111101011", "111011111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "000001000010", "000110010101", "000110010101", "001111001010", "000101000010", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "000001000010", "000001100011", "000001000010", "001111001010", "001111001010", "000001100011", "010001000100", "110111011011", "111011111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "000101000010", "000001100011", "000110010101", "000110010101", "000001000010", "010101010101", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "000001100011", "000110010101", "000001000010", "000110010101", "001111001010", "000110010101", "010101010101", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "000001000010", "000001100011", "000001100011", "000001000010", "010101010101", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "000101100011", "000110010101", "000001100011", "000001000010", "001111001010", "000110010101", "010101010101", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "001000100010", "010100001001", "010100001001", "001000100010", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101100", "010001000100", "000001100011", "000001100011", "000001000010", "000110010101", "001000100010", "010001000100", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "100000111100", "100000111100", "010100001001", "001000000110", "001100000111", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011111110", "010101010101", "001000100010", "100000111100", "010100001001", "001000100010", "010100001001", "011000011001", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011000011001", "001000000110", "001000000110", "000100000011", "000100000011", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "100000111100", "001000000110", "001000000110", "100000111100", "100000111100", "010100001001", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001000100", "100000111100", "010100001001", "001000000110", "001000000110", "001000100010", "110111101100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "001000000011", "010100001001", "100000111100", "010100001001", "010100001001", "001000000110", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "001100000111", "001000000110", "111010101011", "000100000011", "111010101011", "011001100110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011001100110", "001100000111", "010100001001", "001000000110", "001000000110", "010100001001", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101011", "010001000100", "010100001001", "111010101011", "000100000011", "111010101011", "100001000101", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101011", "010001000100", "001000000110", "100000111100", "010100001001", "001000100010", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101011", "010001000100", "111010101011", "101101111000", "000100000011", "101101111000", "111010101011", "010001000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "100000111100", "001000000110", "001000000110", "001000100010", "010101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "101101111000", "111011101110", "001000100010", "010100001001", "001000100010", "111011101110", "101101111000", "011001100110", "111011111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "010001000100", "001000100010", "010100001001", "010100001001", "001000100010", "010001000100", "111011101101", "111111111111", "111111111111", "111111111110", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "111010101011", "111011101110", "001000100010", "010100001001", "001000100010", "111010101011", "111011101110", "101101111000", "010001000100", "011001100110", "011001100110", "011001100110", "011001100110", "010101010101", "011001100110", "011001100110", "010101010101", "010001000100", "001000100010", "001000100010", "100000111100", "001000000110", "001000100010", "001000100010", "010001000100", "011001100110", "011101110111", "011101110111", "011101110111", "100110011001", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110010001001", "111011101110", "101101111000", "001000100010", "000100000011", "001000100010", "101101111000", "111011101110", "111011101110", "001000100010", "101101111000", "111010101011", "111010101011", "111010101011", "111011101110", "111011101110", "111011101110", "111011101110", "111010101011", "111010101011", "001000100010", "100000111100", "001000000110", "001000100010", "101101111000", "111011101110", "111010101011", "001000100010", "101101111000", "111010101011", "101101111000", "011001100110", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101100", "100010001000", "110111101011", "110111101011", "011001100110", "111110111100", "111011101110", "001000100010", "101101111000", "100001000101", "001000100010", "101101111000", "111011101110", "111011101110", "101101111000", "001000100010", "101101111000", "101101111000", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000000110", "000100000011", "100000111100", "001000100010", "001000100010", "101101111000", "101101111000", "001000100010", "101101111000", "101101111000", "100001000101", "011101110111", "111011111110", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "110111101011", "011001100110", "011000101010", "010001000100", "010001000100", "100101001101", "111010101011", "111010101011", "001000100010", "111010101011", "101101111000", "001000100010", "111010101011", "111011101110", "111011101110", "111010101011", "001000100010", "100001000101", "001000100010", "100001000101", "101101111000", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "001000100010", "001000000110", "000100000011", "100000111100", "001000000110", "001000100010", "100001000101", "100001000101", "001000100010", "100001000101", "100001000101", "100001000101", "010101010101", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "010001000100", "001000100010", "001000100010", "010100001001", "001000000110", "101101111000", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "001000100010", "001000100010", "100001000101", "001000100010", "001000100010", "001000100010", "101101111000", "111010101011", "111010101011", "111010101011", "001000100010", "000100000011", "100000111100", "100000111100", "010100001001", "001000100010", "101101111000", "101101111000", "001000100010", "101101111000", "101101111000", "100001000101", "010001000100", "110111101011", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101100", "011001100110", "101101111000", "111010101011", "111010101011", "100001000101", "001000100010", "001000100010", "001000100010", "100001000101", "101101111000", "111010101011", "111010101011", "111010101011", "101101111000", "111010101011", "111010101011", "111010101011", "101101111000", "101101111000", "001000100010", "101101111000", "101101111000", "101101111000", "100001000101", "001000100010", "100001000101", "101101111000", "101101111000", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "001000100010", "011001100110", "110111101011", "111011111110", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "101010101010", "101110001001", "101101111000", "101101111000", "001000100010", "101101111000", "101101111000", "101101111000", "100001000101", "001000100010", "100001000101", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "100001000101", "001000100010", "100001000101", "101101111000", "111010101011", "111010101011", "101101111000", "100001000101", "001000100010", "100001000101", "001000100010", "100001000101", "101101111000", "111010101011", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111010101011", "101101111000", "100001000101", "100001000101", "100001000101", "010001000100", "100010001000", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011001100110", "100001000101", "101101111000", "101101111000", "100001000101", "100001000101", "010001000100", "010101010101", "010101010101", "010001000100", "100001000101", "101101111000", "101101111000", "101101111000", "101101111000", "100001000101", "001000100010", "001000100010", "100001000101", "100001000101", "100001000101", "100001000101", "100001000101", "100001000101", "100001000101", "100001000101", "001000100010", "100001000101", "101101111000", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "111010101011", "101101111000", "101101111000", "100001000101", "100101100111", "111011101110", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011101110111", "011001100110", "011001100110", "011001100110", "011101110111", "110111101100", "111011101101", "111011101101", "110011011011", "010001000100", "101101111000", "101101111000", "101101111000", "100001000101", "010001000100", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010001000100", "100001000101", "100001000101", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "101101111000", "100001000101", "100001000101", "100001000101", "010001000100", "011101110111", "111111111110", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "010101010101", "100001000101", "101101111000", "100001000101", "010001000100", "110011011011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "010101010101", "011101110111", "110111101011", "111011101101", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011101110111", "100001000101", "101101111000", "100001000101", "010101010101", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111101100", "010001000100", "101101111000", "010001000100", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "010101010101", "101101111000", "010101010101", "110111101011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101010110", "011101110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111")

);

begin

row <= GreenGoblin_ROM(conv_integer(address(11 downto 6)));
pixel_out <= row(conv_integer(address(5 downto 0)));

end Behavioral;
