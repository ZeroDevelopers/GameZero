----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 29.04.2017 18:34:01
-- Design Name: 
-- Module Name: player1_rom - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SilverSurfer_4_rom is
    Port ( address : in STD_LOGIC_VECTOR (11 downto 0);
           pixel_out : out STD_LOGIC_VECTOR (11 downto 0));
end SilverSurfer_4_rom;

architecture Behavioral of SilverSurfer_4_rom is

type row_type is array(0 to 63) of std_logic_vector(11 downto 0);
type SilverSurfer_4_rom_type is array(0 to 63) of row_type;
signal row : row_type;

constant SilverSurfer_4_ROM : SilverSurfer_4_rom_type := 
(
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011100", "101110101001", "101110011001", "101110101010", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011101000100", "101001000101", "111010011000", "110001100110", "100001100110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101110", "100101100111", "100001101000", "111010011000", "111011101110", "111011001100", "110001110111", "110010111011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111011100", "101001010110", "001010101101", "110110111100", "111011101110", "111011001100", "101101010110", "110010111010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "101001010110", "001010101101", "110110101010", "111010111010", "111011011100", "110001100101", "101010000111", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "100101110111", "001010011100", "100001111000", "111110000110", "111111011101", "111110000110", "100101100101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "110011011101", "010010001001", "000110111110", "000111001110", "001110011101", "110011011101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110010101010", "011100110101", "011100110101", "110101110101", "110101110110", "111010000110", "101110101001", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "110010101001", "011010010111", "000110111110", "001011101111", "001111111111", "001111111111", "001111101111", "001011001110", "011110111101", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "011000110100", "101001000101", "111010111010", "011101000011", "101101010110", "110010111010", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011100", "101001110110", "010110001000", "001011101111", "010111111111", "011111111111", "001111111111", "001111111111", "010111111111", "011111111111", "001111101111", "010111001101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "111011011101", "110010111010", "101010011000", "100101100110", "100100110100", "101101010101", "111110011000", "110010001000", "100001000100", "100101110111", "100101110111", "101001110111", "100001010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "100101110110", "011001111000", "001011001110", "001111111111", "001111111111", "010011111111", "101111111111", "111011111111", "001111111111", "010011111111", "001111111111", "001111101111", "010010011101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100110000111", "010100100011", "011100100100", "110001010101", "111110000110", "101101010101", "111001110101", "111110000110", "111110000110", "111001110101", "110110011001", "111011011101", "111011001011", "101001010110", "100101100101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110011001011", "101101110110", "010110011010", "001111101111", "110111111111", "011011111111", "111111111111", "111111111111", "111111111111", "111111111111", "100111111111", "101111111111", "001111111111", "010011001101", "110111011101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "101010001000", "101001100111", "110101110110", "111010101001", "111011001100", "110001100101", "101101000101", "111110101001", "111110101000", "110110000111", "110110101010", "111111001011", "111011011101", "111011001011", "110001110111", "011100110100", "100101110110", "100101110111", "101110011001", "111011101110", "110111011101", "101010001000", "100101110110", "100101110110", "110010101001", "111011011101", "110010111011", "100001010100", "010101000100", "001011001110", "001111111111", "001111111111", "100111111111", "111111111111", "111111111111", "111111111111", "111111111111", "101111111111", "010011111111", "001111111111", "001111011111", "100011001110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011000110011", "111001110101", "101001010110", "101011001101", "111111011101", "110001100101", "011001000110", "101011001100", "111111111111", "111111111111", "111011101110", "110110101001", "110110101010", "110110000111", "101000110101", "100100110100", "110001110110", "110010011001", "110001110111", "100101100110", "100101010110", "101001000101", "110001110101", "110001110110", "101001100110", "100101100110", "101101110111", "100000110100", "010101000110", "001011011111", "001111111111", "001111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011011111111", "001111111111", "001111101111", "100011011110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "010100110100", "100101010110", "010100100100", "010110111101", "011110111100", "101001100110", "011001000110", "010110111100", "111011001100", "111011011100", "110110001000", "101001010101", "100101000101", "100000110101", "011100110101", "100000100100", "110001010101", "110110000111", "110101100110", "101001000101", "101001000101", "101101010101", "110110000111", "110110011001", "110010001000", "101001000101", "100100110100", "100000100100", "011000110110", "000110111110", "001111111111", "001111111111", "011111111111", "111111111111", "111111111111", "111111111111", "111111111111", "101011111111", "001111111111", "001111111111", "001011011111", "011110111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "010100110100", "100001100111", "010000100011", "001001101001", "000010111110", "100001100111", "011100110101", "000010101101", "000010111110", "101110000111", "110101110101", "011001010111", "010001101000", "010100110101", "011100110100", "100000110101", "100000100100", "100100110100", "100000110101", "010001101001", "011001000111", "100000100100", "100101000101", "100001000110", "100101000101", "011001010111", "011100110101", "001001111010", "010100110101", "010001111001", "001011101111", "110111111111", "011011111111", "110111111111", "111111111111", "111111111111", "110111111111", "100011111111", "101111111111", "001111111111", "010011001110", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011000110011", "011101010111", "010000110110", "010100100100", "011001010111", "100100100100", "100000100100", "011100110101", "010001111001", "010101011000", "100000100100", "011000100011", "010100110100", "100110001000", "101010001000", "010101000110", "010100110101", "011100100100", "010101000110", "000110001010", "010101000110", "100000110101", "010001011000", "001101111001", "010001101000", "011101101000", "101010011001", "100101010111", "011001000100", "010001101000", "001111001110", "001111111111", "010011111111", "010111111111", "100111111111", "101011111111", "010011111111", "010111111111", "001111111111", "001111101111", "011110101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011000110011", "010101111001", "010000110110", "010100100011", "001001111010", "100101000110", "100100110100", "110001100101", "101101010101", "101101010101", "100000100100", "011100100011", "010000100011", "111111111111", "111111111111", "100110001000", "100110001000", "101010001000", "100110001000", "100110001000", "100101110111", "011000110101", "010000110101", "011101000101", "100110001000", "110010111100", "111111111111", "111011101110", "111111101110", "111111111110", "101111101110", "010011101111", "010011111111", "010111111111", "001111111111", "001111111111", "010011111111", "010111111111", "001011011111", "101011011101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011100", "010100110100", "001010101100", "100100100100", "100000110100", "001001111001", "100110001000", "101001000101", "111010000111", "111111001011", "111011001011", "111010000111", "101101010101", "011000100011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "101110011001", "100110000111", "110010111010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011111111", "001110101110", "001011011111", "001111111111", "001111111111", "001111101111", "000110111110", "100110111100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100110000111", "011101000110", "000110011100", "100100100100", "100100110100", "010000100011", "001001111010", "111001110110", "111001110101", "111111101110", "111011011100", "111010011000", "100100110100", "011100100100", "010000100010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "011110101100", "001010111110", "001111001110", "010110101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "100101110111", "101001010110", "100101000110", "101101000101", "100001010101", "110111001011", "100001110111", "001101101000", "100101000110", "110110000111", "111011001011", "110001010101", "100000100100", "101001000101", "011000100011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "100001000101", "001001111010", "101001000101", "100000110100", "110111001011", "111111111111", "111111111110", "011000110100", "100000100100", "110001100110", "111010111010", "111001110101", "100100110100", "100000100100", "011101000100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "100001000101", "000110101101", "100000100100", "010100100011", "110111001100", "111111111111", "111011101101", "011000110011", "101001000101", "111001110101", "111010101001", "110101110111", "110101100101", "100100110100", "100001010101", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "011001000100", "001101111010", "100000100100", "101101010101", "110010111010", "111111111111", "100101110111", "101001000101", "111110000110", "111010101001", "111011101110", "111011101110", "111110010111", "111001110101", "100101100110", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "100101110111", "101001000101", "011000110101", "111010010111", "101110001000", "111111111111", "101010001000", "110110011000", "111110011000", "100010111100", "111011101110", "111111101110", "111110111001", "111001110101", "101001000101", "100001010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "000110101101", "010100110110", "111110101001", "101010001000", "111111111111", "100110001000", "111010111010", "111110011000", "001111001110", "111011101110", "111011001011", "111010101001", "111110000110", "110001100101", "011100100100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "101010001000", "001110001010", "011101000110", "111110010111", "101001110111", "111111111111", "100001010110", "001010101101", "110010111010", "100101010110", "010110111101", "011010111100", "000110111110", "110101100101", "111001110101", "101001000101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "010000110100", "011001000111", "111001110101", "100001000101", "110010111010", "100000110101", "001101000111", "000010101101", "011100100100", "001001101001", "000010111110", "000110011011", "110001010101", "111110101000", "101101010101", "100001010100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011001010101", "001101011000", "100000100100", "011000100011", "100101000101", "010100110101", "100000100100", "011001000110", "100000100100", "011000100100", "010101000111", "011100100100", "110001100110", "111010111010", "111001110110", "100001010110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111011100", "010001111010", "101001000101", "100000110100", "010000100011", "000110011100", "001001111010", "100000100100", "011100100100", "010000100011", "001101011000", "011001000110", "110001010101", "111010111010", "111010111010", "100101010101", "101110011001", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "010010001010", "011100110011", "011000100011", "001100110100", "000010111110", "000010101101", "011100110101", "011101000101", "011100110011", "000010101101", "011001010111", "100100110100", "111010011000", "111111111111", "110001110111", "100001100110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "010001111001", "010000100011", "010000100100", "001101011000", "000011001111", "000010101101", "011100110101", "110001010101", "011100110011", "100001100111", "011001010111", "100100110100", "111010000111", "111111111111", "111110111001", "100001100110", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "100001111000", "010001011000", "010100100011", "001001111010", "000011001111", "000110101101", "100100110101", "111110000101", "011100110011", "010101000101", "100001111000", "100000100100", "110101100101", "111011011101", "111011011101", "100001100110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "011101010101", "010100100011", "000011001111", "000011001111", "010000110110", "101001000101", "111001110101", "011000110100", "010101000101", "000010101101", "100000100100", "110101100101", "111110111010", "111111111111", "011100110100", "011101010101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "100001110110", "000011001111", "000110001011", "011100110101", "110101110101", "110001100101", "110010111010", "110111001100", "001110011011", "011001101000", "100100110100", "111110000110", "111111101110", "100000110101", "101110101000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "000110111110", "011001000110", "101001000100", "111110000110", "100000110101", "111111111111", "111111111111", "100101110111", "010001111010", "100100110101", "110001010101", "111011001011", "101001010110", "110010111010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "100101110110", "100001100111", "011000110101", "110101100101", "101101010101", "100001100110", "111111111111", "111111111111", "110111001011", "011001010111", "011100110101", "100100110100", "111110000110", "101001010101", "110010111011", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111011100", "101001010110", "101001000101", "010001101000", "100000100100", "100001010110", "111111101110", "111111111111", "111111111111", "111111111111", "110111001100", "100000110101", "100000100100", "110001010101", "100000110101", "110010101001", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "100101110111", "100101000101", "011100110101", "011000110101", "100000110101", "101110101001", "111111111111", "111111111111", "111111111111", "111111111111", "111011101110", "010101000111", "010001011000", "101001000101", "100000100100", "011101000101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111001100", "011001000101", "101001010110", "100000100100", "100000100100", "100000110101", "111011011101", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "010101000111", "001101101001", "100000100100", "101001000110", "100001100110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111001100", "011010001001", "000010111110", "011101111000", "100000100100", "100000110101", "100001110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111001100", "010101000110", "010100110110", "100000100100", "110001100110", "100001100110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "010101000101", "000110011100", "000010111110", "011101101000", "100100110100", "100001010101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "011001000101", "000110101101", "010100110110", "100000100100", "101101010101", "101010011000", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "101110101001", "011000110101", "000010101101", "001010011011", "100000110101", "101101010101", "101010001000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "010001010110", "000010111110", "100100110100", "110101110110", "011000110100", "100001110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100110000111", "101101010101", "011001101000", "101001000101", "101001000101", "100000110101", "110010111010", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "010001010110", "000010111110", "101000110100", "111010111011", "001100100010", "100001110111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "101101010101", "101101010101", "100000100100", "100100110101", "100001100110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "011001000101", "001010001011", "100100110100", "111111011100", "010101010101", "100110000111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "100001100111", "100001100111", "100000100100", "011101000101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "100001010110", "101001000101", "101001000101", "111010101001", "011101010101", "100101100111", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "001010001011", "100001100111", "100000100100", "101110011001", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011100", "100001010110", "010101111001", "101001000101", "011001000011", "011101000101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "010101111001", "101101000101", "100000110101", "110111011100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "101010001000", "011001010111", "100001000110", "111001110101", "011101000101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "101101010101", "010101111001", "011101000100", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "011101010101", "011101111000", "100000100100", "011101000100", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "101101000101", "001110001010", "011101000101", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110010111010", "100001010111", "100000100100", "011101000100", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "100101110111", "101101010101", "100001000110", "011001000100", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "110111001011", "001110001010", "100000100100", "011101000100", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "111111111111", "111111111111", "111111101110", "100001100110", "101101000101", "100100110100", "001010001011", "110010111011", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101101", "101110011001", "001010101100", "100100100100", "011101000100", "111011011100", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "111011011100", "100101110111", "100110000111", "100101110111", "100101010110", "100000110101", "100000110101", "100000110101", "011000100011", "101001000101", "100100110100", "010101000110", "011100110100", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "011000110011", "101001010101", "100100110100", "100101000101", "100001100110", "111011101110", "111111101110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101110", "011101010101", "011101000100", "010101000101", "011101000110", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "100101000100", "011101000101", "000110111101", "101001010101", "100000100100", "011000100011", "100101000100", "100101000100", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101001000101", "011000100011", "101001000101", "100000100100", "110010001000", "011100100100", "011100110100", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100000110101", "100001010101", "100001100110", "100001110110", "100001110110", "100110001000", "111111111111", "111111111111"), 
("011000110100", "100001010110", "110111001100", "111011011101", "111111111111", "101110001000", "001101111001", "001010101100", "000010111110", "000010101101", "100110011001", "111010000111", "111001110101", "111001110101", "111001110101", "010100100010", "010001101001", "000010111110", "100001100111", "100000100100", "100100110101", "011100100100", "100101000100", "011100110011", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "011100110011", "100101010110", "100101010110", "101001000101", "110001010101", "011100100100", "010100100011", "101001000101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "101101010101", "100100110101", "100100110101", "100001010110", "011101000100"), 
("110010011001", "110110001000", "101001010101", "101001100111", "111111111111", "100000100100", "101101010101", "001101111010", "001010101100", "001110111101", "000010111110", "000011001111", "000011001111", "101110101010", "101110011000", "010001000101", "010100110101", "001101101000", "100000110100", "011100100100", "011100100100", "100101000100", "100000110100", "100001000011", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "011100110011", "100001100111", "000110101101", "011001101000", "100100100100", "101101010110", "110101110110", "011100100011", "110001100101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "111001110101", "110101110110"), 
("110010000111", "100000110100", "010000100010", "100001100110", "111111111111", "011001000100", "010100110011", "010100100011", "011000100011", "100101000101", "011101010111", "011101111000", "000110011100", "000110011100", "000010111110", "000010111110", "000110011011", "000110011011", "000110011011", "000110011011", "000110011011", "000110011011", "000110011011", "010010111100", "010010111100", "010010111100", "010010111100", "010010111100", "010010111100", "010010111100", "001010011100", "010100100100", "000011001111", "001010101100", "100100110100", "101101010110", "111010111010", "101101010101", "010100100011", "011001000100", "101101100101", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110000110", "111110010111", "111110101000", "111110111010", "111011011101", "111111011101", "110110111011"), 
("010100100011", "010100110011", "011001000100", "110010111011", "111111111111", "111011101101", "101110101001", "100001100110", "010100100011", "010000100010", "010000100010", "010000100010", "011000100011", "011100100100", "011100100100", "100101000100", "010101010111", "001001101001", "001001101001", "000110011100", "001010011100", "001010011100", "001010101100", "001010101100", "001010101100", "001010101100", "001010101100", "001010101100", "001010101100", "001010101100", "001010101100", "001110001010", "011101100111", "100001010111", "011000100011", "010100100011", "011000110011", "011001010111", "010001000110", "101101100110", "010100100011", "111010111010", "111010111010", "111010111010", "111010111010", "111010111010", "111010111010", "111010111010", "111111011100", "111111011100", "111111011100", "111111011100", "111111011100", "111111011100", "111111011100", "111111011100", "111111011101", "111011011100", "111010111010", "111110101000", "110001111000", "101001010110", "011100110011", "011000100011"), 
("100001100110", "101110101001", "111011101101", "111111111111", "111111111111", "111111111111", "111111111111", "111011011101", "001110001001", "100101000100", "100000110100", "011100100100", "011100100100", "011100100100", "010100110011", "011001000100", "011001000100", "010100110100", "010100110011", "010100100011", "010100100011", "010100100011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000100011", "011000100011", "001110001010", "001010101100", "001010101100", "011000100011", "011000100011", "011000100011", "110010101010", "111011001100", "111011001100", "111011001100", "111011001100", "111011001100", "111011001100", "111011001100", "110111001100", "110110101010", "110110001000", "110010000111", "110001110101", "110001100101", "101001000100", "100101000100", "100101000100", "011100100100", "011100100100", "010000100011", "010100110011", "010100110011", "010100110011", "011101010101"), 
("111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "001110101011", "101101010101", "100101010111", "100101000101", "011000110100", "100001100110", "110111001100", "111111111111", "111111111111", "111111111111", "101110011001", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000110011", "011000100011", "010100100011", "010100100011", "010000100010", "010000100010", "010000100010", "010000100010", "010100100011", "010100110100", "011000110100", "011001000100", "100101110111", "110010111010", "110010111011", "110111001011", "111011101101"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "001110101011", "101001010110", "001101101001", "010100110100", "101010001000", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100001100110", "100101110111", "110111011100", "111011101101", "111111101110", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111110", "010110011011", "010001111010", "011101010110", "100101110111", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111101110", "111111111110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111011101101", "111011011101", "111111101110", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"), 
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111"),
("111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111", "111111111111")

);

begin

row <= SilverSurfer_4_ROM(conv_integer(address(11 downto 6)));
pixel_out <= row(conv_integer(address(5 downto 0)));

end Behavioral;